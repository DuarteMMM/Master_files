VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO test
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN test 0 0 ;
  SIZE 28.5 BY 85 ;
  SYMMETRY X Y R90 ;
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME3 ;
        RECT 14.2 84 15.2 85 ;
    END
  END dvdd
  PIN cc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 19.3 28.5 20.3 ;
    END
  END cc
  PIN tc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 17.8 28.5 18.8 ;
    END
  END tc
  PIN cv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 16.3 28.5 17.3 ;
    END
  END cv
  PIN imonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 14.8 28.5 15.8 ;
    END
  END imonen
  PIN vmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 13.3 28.5 14.3 ;
    END
  END vmonen
  PIN tmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 11.8 28.5 12.8 ;
    END
  END tmonen
  PIN vtok
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 8.5 0 9.5 1 ;
    END
  END vtok
  PIN ibat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 59.8 1 60.8 ;
    END
  END ibat[7]
  PIN ibat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 49.3 1 50.3 ;
    END
  END ibat[0]
  PIN tbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 47.3 1 48.3 ;
    END
  END tbat[7]
  PIN vcutoff[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 24.3 1 25.3 ;
    END
  END vcutoff[0]
  PIN vpreset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 11.8 1 12.8 ;
    END
  END vpreset[0]
  PIN tempmin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 72.3 28.5 73.3 ;
    END
  END tempmin[7]
  PIN tempmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 50.8 28.5 51.8 ;
    END
  END tempmax[1]
  PIN tempmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 49.3 28.5 50.3 ;
    END
  END tempmax[0]
  PIN iend[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 34.8 28.5 35.8 ;
    END
  END iend[7]
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME3 ;
        RECT 10 0 11 1 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 11.5 0 12.5 1 ;
    END
  END en
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 14.5 0 15.5 1 ;
    END
  END rstz
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 17.5 0 18.5 1 ;
    END
  END si
  PIN se
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 16 0 17 1 ;
    END
  END se
  PIN so
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 19 0 20 1 ;
    END
  END so
  PIN ibat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 50.8 1 51.8 ;
    END
  END ibat[1]
  PIN tbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 36.8 1 37.8 ;
    END
  END tbat[0]
  PIN ibat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 52.3 1 53.3 ;
    END
  END ibat[2]
  PIN ibat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 53.8 1 54.8 ;
    END
  END ibat[3]
  PIN ibat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 55.3 1 56.3 ;
    END
  END ibat[4]
  PIN ibat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 56.8 1 57.8 ;
    END
  END ibat[5]
  PIN ibat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 58.3 1 59.3 ;
    END
  END ibat[6]
  PIN vbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 61.8 1 62.8 ;
    END
  END vbat[0]
  PIN vbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 72.3 1 73.3 ;
    END
  END vbat[7]
  PIN vbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 63.3 1 64.3 ;
    END
  END vbat[1]
  PIN vbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 64.8 1 65.8 ;
    END
  END vbat[2]
  PIN vbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 66.3 1 67.3 ;
    END
  END vbat[3]
  PIN vbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 67.8 1 68.8 ;
    END
  END vbat[4]
  PIN vbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 69.3 1 70.3 ;
    END
  END vbat[5]
  PIN vbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 70.8 1 71.8 ;
    END
  END vbat[6]
  PIN tbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 38.3 1 39.3 ;
    END
  END tbat[1]
  PIN tbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 45.8 1 46.8 ;
    END
  END tbat[6]
  PIN tbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 41.3 1 42.3 ;
    END
  END tbat[3]
  PIN tbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 44.3 1 45.3 ;
    END
  END tbat[5]
  PIN tbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 42.8 1 43.8 ;
    END
  END tbat[4]
  PIN tbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 39.8 1 40.8 ;
    END
  END tbat[2]
  PIN vcutoff[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 28.8 1 29.8 ;
    END
  END vcutoff[3]
  PIN vcutoff[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 34.8 1 35.8 ;
    END
  END vcutoff[7]
  PIN vcutoff[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 25.8 1 26.8 ;
    END
  END vcutoff[1]
  PIN vcutoff[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 27.3 1 28.3 ;
    END
  END vcutoff[2]
  PIN vcutoff[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 30.3 1 31.3 ;
    END
  END vcutoff[4]
  PIN vcutoff[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 33.3 1 34.3 ;
    END
  END vcutoff[6]
  PIN vcutoff[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 31.8 1 32.8 ;
    END
  END vcutoff[5]
  PIN tempmin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 66.3 28.5 67.3 ;
    END
  END tempmin[3]
  PIN tempmin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 63.3 28.5 64.3 ;
    END
  END tempmin[1]
  PIN tempmin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 67.8 28.5 68.8 ;
    END
  END tempmin[4]
  PIN tempmin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 70.8 28.5 71.8 ;
    END
  END tempmin[6]
  PIN tempmin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 64.8 28.5 65.8 ;
    END
  END tempmin[2]
  PIN tempmin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 69.3 28.5 70.3 ;
    END
  END tempmin[5]
  PIN tempmin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 61.8 28.5 62.8 ;
    END
  END tempmin[0]
  PIN vpreset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 19.3 1 20.3 ;
    END
  END vpreset[5]
  PIN vpreset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 14.8 1 15.8 ;
    END
  END vpreset[2]
  PIN vpreset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 20.8 1 21.8 ;
    END
  END vpreset[6]
  PIN vpreset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 17.8 1 18.8 ;
    END
  END vpreset[4]
  PIN vpreset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 13.3 1 14.3 ;
    END
  END vpreset[1]
  PIN vpreset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 16.3 1 17.3 ;
    END
  END vpreset[3]
  PIN vpreset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 0 22.3 1 23.3 ;
    END
  END vpreset[7]
  PIN tempmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 52.3 28.5 53.3 ;
    END
  END tempmax[2]
  PIN tempmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 59.8 28.5 60.8 ;
    END
  END tempmax[7]
  PIN tempmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 58.3 28.5 59.3 ;
    END
  END tempmax[6]
  PIN tempmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 56.8 28.5 57.8 ;
    END
  END tempmax[5]
  PIN tempmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 55.3 28.5 56.3 ;
    END
  END tempmax[4]
  PIN tempmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 53.8 28.5 54.8 ;
    END
  END tempmax[3]
  PIN tmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 36.8 28.5 37.8 ;
    END
  END tmax[0]
  PIN tmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 39.8 28.5 40.8 ;
    END
  END tmax[2]
  PIN tmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 38.3 28.5 39.3 ;
    END
  END tmax[1]
  PIN tmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 41.3 28.5 42.3 ;
    END
  END tmax[3]
  PIN tmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 42.8 28.5 43.8 ;
    END
  END tmax[4]
  PIN tmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 44.3 28.5 45.3 ;
    END
  END tmax[5]
  PIN tmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 45.8 28.5 46.8 ;
    END
  END tmax[6]
  PIN tmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 47.3 28.5 48.3 ;
    END
  END tmax[7]
  PIN iend[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 33.3 28.5 34.3 ;
    END
  END iend[6]
  PIN iend[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 31.8 28.5 32.8 ;
    END
  END iend[5]
  PIN iend[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 30.3 28.5 31.3 ;
    END
  END iend[4]
  PIN iend[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 28.8 28.5 29.8 ;
    END
  END iend[3]
  PIN iend[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 27.3 28.5 28.3 ;
    END
  END iend[2]
  PIN iend[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 25.8 28.5 26.8 ;
    END
  END iend[1]
  PIN iend[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 27.5 24.3 28.5 25.3 ;
    END
  END iend[0]
  PIN dgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME3 ;
        RECT 13 0 14 1 ;
    END
  END dgnd
  OBS
    LAYER ME1 SPACING 0.16 ;
      RECT 0 0 28.5 85 ;
    LAYER ME2 SPACING 0.2 ;
      RECT 0 0 28.5 85 ;
    LAYER ME3 SPACING 0.2 ;
      RECT 15.56 73.66 28.5 85 ;
      RECT 0 73.66 13.84 85 ;
      RECT 1.36 1.36 27.14 83.64 ;
      RECT 0 61.16 28.5 61.44 ;
      RECT 0 48.66 28.5 48.94 ;
      RECT 0 36.16 28.5 36.44 ;
      RECT 0 23.66 28.5 23.94 ;
      RECT 1.36 20.66 28.5 23.94 ;
      RECT 20.36 0 28.5 11.44 ;
      RECT 0 0 8.14 11.44 ;
    LAYER ME4 SPACING 0.2 ;
      RECT 15.5 73.6 28.5 85 ;
      RECT 0 73.6 13.9 85 ;
      RECT 1.3 1.3 27.2 83.7 ;
      RECT 0 61.1 28.5 61.5 ;
      RECT 0 48.6 28.5 49 ;
      RECT 0 36.1 28.5 36.5 ;
      RECT 0 23.6 28.5 24 ;
      RECT 1.3 20.6 28.5 24 ;
      RECT 20.3 0 28.5 11.5 ;
      RECT 0 0 8.2 11.5 ;
    LAYER ME5 SPACING 0.2 ;
      RECT 0 0 28.5 85 ;
    LAYER ME6 SPACING 0.2 ;
      RECT 0 0 28.5 85 ;
    LAYER ME7 SPACING 0.4 ;
      RECT 0 0 28.5 85 ;
    LAYER ME8 SPACING 1.5 ;
      RECT 0 0 28.5 85 ;
  END
END test

END LIBRARY
