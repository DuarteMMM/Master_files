##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Sun Jan  8 15:21:40 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERctr
  CLASS BLOCK ;
  SIZE 47.200000 BY 68.000000 ;
  FOREIGN BATCHARGERctr 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN cc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 26.100000 0.520000 26.300000 ;
    END
  END cc
  PIN tc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 28.100000 0.520000 28.300000 ;
    END
  END tc
  PIN cv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 30.100000 0.520000 30.300000 ;
    END
  END cv
  PIN imonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 32.100000 0.520000 32.300000 ;
    END
  END imonen
  PIN vmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 34.100000 0.520000 34.300000 ;
    END
  END vmonen
  PIN tmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 36.100000 0.520000 36.300000 ;
    END
  END tmonen
  PIN vtok
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 20.100000 0.520000 20.300000 ;
    END
  END vtok
  PIN vbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 5.700000 47.200000 5.900000 ;
    END
  END vbat[7]
  PIN vbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 4.900000 47.200000 5.100000 ;
    END
  END vbat[6]
  PIN vbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 4.100000 47.200000 4.300000 ;
    END
  END vbat[5]
  PIN vbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 3.300000 47.200000 3.500000 ;
    END
  END vbat[4]
  PIN vbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 2.500000 47.200000 2.700000 ;
    END
  END vbat[3]
  PIN vbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 1.700000 47.200000 1.900000 ;
    END
  END vbat[2]
  PIN vbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 0.900000 47.200000 1.100000 ;
    END
  END vbat[1]
  PIN vbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 0.100000 47.200000 0.300000 ;
    END
  END vbat[0]
  PIN ibat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 12.500000 47.200000 12.700000 ;
    END
  END ibat[7]
  PIN ibat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 11.700000 47.200000 11.900000 ;
    END
  END ibat[6]
  PIN ibat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 10.900000 47.200000 11.100000 ;
    END
  END ibat[5]
  PIN ibat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 10.100000 47.200000 10.300000 ;
    END
  END ibat[4]
  PIN ibat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 9.300000 47.200000 9.500000 ;
    END
  END ibat[3]
  PIN ibat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 8.500000 47.200000 8.700000 ;
    END
  END ibat[2]
  PIN ibat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 7.700000 47.200000 7.900000 ;
    END
  END ibat[1]
  PIN ibat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 6.900000 47.200000 7.100000 ;
    END
  END ibat[0]
  PIN tbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 19.300000 47.200000 19.500000 ;
    END
  END tbat[7]
  PIN tbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 18.500000 47.200000 18.700000 ;
    END
  END tbat[6]
  PIN tbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 17.700000 47.200000 17.900000 ;
    END
  END tbat[5]
  PIN tbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 16.900000 47.200000 17.100000 ;
    END
  END tbat[4]
  PIN tbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 16.100000 47.200000 16.300000 ;
    END
  END tbat[3]
  PIN tbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 15.300000 47.200000 15.500000 ;
    END
  END tbat[2]
  PIN tbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 14.500000 47.200000 14.700000 ;
    END
  END tbat[1]
  PIN tbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 13.700000 47.200000 13.900000 ;
    END
  END tbat[0]
  PIN vcutoff[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 26.100000 47.200000 26.300000 ;
    END
  END vcutoff[7]
  PIN vcutoff[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 25.300000 47.200000 25.500000 ;
    END
  END vcutoff[6]
  PIN vcutoff[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 24.500000 47.200000 24.700000 ;
    END
  END vcutoff[5]
  PIN vcutoff[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 23.700000 47.200000 23.900000 ;
    END
  END vcutoff[4]
  PIN vcutoff[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 22.900000 47.200000 23.100000 ;
    END
  END vcutoff[3]
  PIN vcutoff[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 22.100000 47.200000 22.300000 ;
    END
  END vcutoff[2]
  PIN vcutoff[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 21.300000 47.200000 21.500000 ;
    END
  END vcutoff[1]
  PIN vcutoff[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 20.500000 47.200000 20.700000 ;
    END
  END vcutoff[0]
  PIN vpreset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 32.900000 47.200000 33.100000 ;
    END
  END vpreset[7]
  PIN vpreset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 32.100000 47.200000 32.300000 ;
    END
  END vpreset[6]
  PIN vpreset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 31.300000 47.200000 31.500000 ;
    END
  END vpreset[5]
  PIN vpreset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 30.500000 47.200000 30.700000 ;
    END
  END vpreset[4]
  PIN vpreset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 29.700000 47.200000 29.900000 ;
    END
  END vpreset[3]
  PIN vpreset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 28.900000 47.200000 29.100000 ;
    END
  END vpreset[2]
  PIN vpreset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 28.100000 47.200000 28.300000 ;
    END
  END vpreset[1]
  PIN vpreset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 27.300000 47.200000 27.500000 ;
    END
  END vpreset[0]
  PIN tempmin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 39.700000 47.200000 39.900000 ;
    END
  END tempmin[7]
  PIN tempmin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 38.900000 47.200000 39.100000 ;
    END
  END tempmin[6]
  PIN tempmin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 38.100000 47.200000 38.300000 ;
    END
  END tempmin[5]
  PIN tempmin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 37.300000 47.200000 37.500000 ;
    END
  END tempmin[4]
  PIN tempmin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 36.500000 47.200000 36.700000 ;
    END
  END tempmin[3]
  PIN tempmin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 35.700000 47.200000 35.900000 ;
    END
  END tempmin[2]
  PIN tempmin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 34.900000 47.200000 35.100000 ;
    END
  END tempmin[1]
  PIN tempmin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 34.100000 47.200000 34.300000 ;
    END
  END tempmin[0]
  PIN tempmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 46.500000 47.200000 46.700000 ;
    END
  END tempmax[7]
  PIN tempmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 45.700000 47.200000 45.900000 ;
    END
  END tempmax[6]
  PIN tempmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 44.900000 47.200000 45.100000 ;
    END
  END tempmax[5]
  PIN tempmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 44.100000 47.200000 44.300000 ;
    END
  END tempmax[4]
  PIN tempmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 43.300000 47.200000 43.500000 ;
    END
  END tempmax[3]
  PIN tempmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 42.500000 47.200000 42.700000 ;
    END
  END tempmax[2]
  PIN tempmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 41.700000 47.200000 41.900000 ;
    END
  END tempmax[1]
  PIN tempmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 40.900000 47.200000 41.100000 ;
    END
  END tempmax[0]
  PIN tmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 53.300000 47.200000 53.500000 ;
    END
  END tmax[7]
  PIN tmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 52.500000 47.200000 52.700000 ;
    END
  END tmax[6]
  PIN tmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 51.700000 47.200000 51.900000 ;
    END
  END tmax[5]
  PIN tmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 50.900000 47.200000 51.100000 ;
    END
  END tmax[4]
  PIN tmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 50.100000 47.200000 50.300000 ;
    END
  END tmax[3]
  PIN tmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 49.300000 47.200000 49.500000 ;
    END
  END tmax[2]
  PIN tmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 48.500000 47.200000 48.700000 ;
    END
  END tmax[1]
  PIN tmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 47.700000 47.200000 47.900000 ;
    END
  END tmax[0]
  PIN iend[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 60.100000 47.200000 60.300000 ;
    END
  END iend[7]
  PIN iend[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 59.300000 47.200000 59.500000 ;
    END
  END iend[6]
  PIN iend[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 58.500000 47.200000 58.700000 ;
    END
  END iend[5]
  PIN iend[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 57.700000 47.200000 57.900000 ;
    END
  END iend[4]
  PIN iend[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 56.900000 47.200000 57.100000 ;
    END
  END iend[3]
  PIN iend[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 56.100000 47.200000 56.300000 ;
    END
  END iend[2]
  PIN iend[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 55.300000 47.200000 55.500000 ;
    END
  END iend[1]
  PIN iend[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.680000 54.500000 47.200000 54.700000 ;
    END
  END iend[0]
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal4 ;
        RECT 23.700000 0.000000 23.900000 0.520000 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 22.100000 0.520000 22.300000 ;
    END
  END en
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 24.100000 0.520000 24.300000 ;
    END
  END rstz
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
        RECT 24.100000 67.480000 24.300000 68.000000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
        RECT 20.100000 67.480000 20.300000 68.000000 ;
    END
  END dgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
    LAYER metal3 ;
      RECT 0.000000 60.500000 47.200000 68.000000 ;
      RECT 0.000000 59.900000 46.480000 60.500000 ;
      RECT 0.000000 59.700000 47.200000 59.900000 ;
      RECT 0.000000 59.100000 46.480000 59.700000 ;
      RECT 0.000000 58.900000 47.200000 59.100000 ;
      RECT 0.000000 58.300000 46.480000 58.900000 ;
      RECT 0.000000 58.100000 47.200000 58.300000 ;
      RECT 0.000000 57.500000 46.480000 58.100000 ;
      RECT 0.000000 57.300000 47.200000 57.500000 ;
      RECT 0.000000 56.700000 46.480000 57.300000 ;
      RECT 0.000000 56.500000 47.200000 56.700000 ;
      RECT 0.000000 55.900000 46.480000 56.500000 ;
      RECT 0.000000 55.700000 47.200000 55.900000 ;
      RECT 0.000000 55.100000 46.480000 55.700000 ;
      RECT 0.000000 54.900000 47.200000 55.100000 ;
      RECT 0.000000 54.300000 46.480000 54.900000 ;
      RECT 0.000000 53.700000 47.200000 54.300000 ;
      RECT 0.000000 53.100000 46.480000 53.700000 ;
      RECT 0.000000 52.900000 47.200000 53.100000 ;
      RECT 0.000000 52.300000 46.480000 52.900000 ;
      RECT 0.000000 52.100000 47.200000 52.300000 ;
      RECT 0.000000 51.500000 46.480000 52.100000 ;
      RECT 0.000000 51.300000 47.200000 51.500000 ;
      RECT 0.000000 50.700000 46.480000 51.300000 ;
      RECT 0.000000 50.500000 47.200000 50.700000 ;
      RECT 0.000000 49.900000 46.480000 50.500000 ;
      RECT 0.000000 49.700000 47.200000 49.900000 ;
      RECT 0.000000 49.100000 46.480000 49.700000 ;
      RECT 0.000000 48.900000 47.200000 49.100000 ;
      RECT 0.000000 48.300000 46.480000 48.900000 ;
      RECT 0.000000 48.100000 47.200000 48.300000 ;
      RECT 0.000000 47.500000 46.480000 48.100000 ;
      RECT 0.000000 46.900000 47.200000 47.500000 ;
      RECT 0.000000 46.300000 46.480000 46.900000 ;
      RECT 0.000000 46.100000 47.200000 46.300000 ;
      RECT 0.000000 45.500000 46.480000 46.100000 ;
      RECT 0.000000 45.300000 47.200000 45.500000 ;
      RECT 0.000000 44.700000 46.480000 45.300000 ;
      RECT 0.000000 44.500000 47.200000 44.700000 ;
      RECT 0.000000 43.900000 46.480000 44.500000 ;
      RECT 0.000000 43.700000 47.200000 43.900000 ;
      RECT 0.000000 43.100000 46.480000 43.700000 ;
      RECT 0.000000 42.900000 47.200000 43.100000 ;
      RECT 0.000000 42.300000 46.480000 42.900000 ;
      RECT 0.000000 42.100000 47.200000 42.300000 ;
      RECT 0.000000 41.500000 46.480000 42.100000 ;
      RECT 0.000000 41.300000 47.200000 41.500000 ;
      RECT 0.000000 40.700000 46.480000 41.300000 ;
      RECT 0.000000 40.100000 47.200000 40.700000 ;
      RECT 0.000000 39.500000 46.480000 40.100000 ;
      RECT 0.000000 39.300000 47.200000 39.500000 ;
      RECT 0.000000 38.700000 46.480000 39.300000 ;
      RECT 0.000000 38.500000 47.200000 38.700000 ;
      RECT 0.000000 37.900000 46.480000 38.500000 ;
      RECT 0.000000 37.700000 47.200000 37.900000 ;
      RECT 0.000000 37.100000 46.480000 37.700000 ;
      RECT 0.000000 36.900000 47.200000 37.100000 ;
      RECT 0.000000 36.500000 46.480000 36.900000 ;
      RECT 0.720000 36.300000 46.480000 36.500000 ;
      RECT 0.720000 36.100000 47.200000 36.300000 ;
      RECT 0.720000 35.900000 46.480000 36.100000 ;
      RECT 0.000000 35.500000 46.480000 35.900000 ;
      RECT 0.000000 35.300000 47.200000 35.500000 ;
      RECT 0.000000 34.700000 46.480000 35.300000 ;
      RECT 0.000000 34.500000 47.200000 34.700000 ;
      RECT 0.720000 33.900000 46.480000 34.500000 ;
      RECT 0.000000 33.300000 47.200000 33.900000 ;
      RECT 0.000000 32.700000 46.480000 33.300000 ;
      RECT 0.000000 32.500000 47.200000 32.700000 ;
      RECT 0.720000 31.900000 46.480000 32.500000 ;
      RECT 0.000000 31.700000 47.200000 31.900000 ;
      RECT 0.000000 31.100000 46.480000 31.700000 ;
      RECT 0.000000 30.900000 47.200000 31.100000 ;
      RECT 0.000000 30.500000 46.480000 30.900000 ;
      RECT 0.720000 30.300000 46.480000 30.500000 ;
      RECT 0.720000 30.100000 47.200000 30.300000 ;
      RECT 0.720000 29.900000 46.480000 30.100000 ;
      RECT 0.000000 29.500000 46.480000 29.900000 ;
      RECT 0.000000 29.300000 47.200000 29.500000 ;
      RECT 0.000000 28.700000 46.480000 29.300000 ;
      RECT 0.000000 28.500000 47.200000 28.700000 ;
      RECT 0.720000 27.900000 46.480000 28.500000 ;
      RECT 0.000000 27.700000 47.200000 27.900000 ;
      RECT 0.000000 27.100000 46.480000 27.700000 ;
      RECT 0.000000 26.500000 47.200000 27.100000 ;
      RECT 0.720000 25.900000 46.480000 26.500000 ;
      RECT 0.000000 25.700000 47.200000 25.900000 ;
      RECT 0.000000 25.100000 46.480000 25.700000 ;
      RECT 0.000000 24.900000 47.200000 25.100000 ;
      RECT 0.000000 24.500000 46.480000 24.900000 ;
      RECT 0.720000 24.300000 46.480000 24.500000 ;
      RECT 0.720000 24.100000 47.200000 24.300000 ;
      RECT 0.720000 23.900000 46.480000 24.100000 ;
      RECT 0.000000 23.500000 46.480000 23.900000 ;
      RECT 0.000000 23.300000 47.200000 23.500000 ;
      RECT 0.000000 22.700000 46.480000 23.300000 ;
      RECT 0.000000 22.500000 47.200000 22.700000 ;
      RECT 0.720000 21.900000 46.480000 22.500000 ;
      RECT 0.000000 21.700000 47.200000 21.900000 ;
      RECT 0.000000 21.100000 46.480000 21.700000 ;
      RECT 0.000000 20.900000 47.200000 21.100000 ;
      RECT 0.000000 20.500000 46.480000 20.900000 ;
      RECT 0.720000 20.300000 46.480000 20.500000 ;
      RECT 0.720000 19.900000 47.200000 20.300000 ;
      RECT 0.000000 19.700000 47.200000 19.900000 ;
      RECT 0.000000 19.100000 46.480000 19.700000 ;
      RECT 0.000000 18.900000 47.200000 19.100000 ;
      RECT 0.000000 18.300000 46.480000 18.900000 ;
      RECT 0.000000 18.100000 47.200000 18.300000 ;
      RECT 0.000000 17.500000 46.480000 18.100000 ;
      RECT 0.000000 17.300000 47.200000 17.500000 ;
      RECT 0.000000 16.700000 46.480000 17.300000 ;
      RECT 0.000000 16.500000 47.200000 16.700000 ;
      RECT 0.000000 15.900000 46.480000 16.500000 ;
      RECT 0.000000 15.700000 47.200000 15.900000 ;
      RECT 0.000000 15.100000 46.480000 15.700000 ;
      RECT 0.000000 14.900000 47.200000 15.100000 ;
      RECT 0.000000 14.300000 46.480000 14.900000 ;
      RECT 0.000000 14.100000 47.200000 14.300000 ;
      RECT 0.000000 13.500000 46.480000 14.100000 ;
      RECT 0.000000 12.900000 47.200000 13.500000 ;
      RECT 0.000000 12.300000 46.480000 12.900000 ;
      RECT 0.000000 12.100000 47.200000 12.300000 ;
      RECT 0.000000 11.500000 46.480000 12.100000 ;
      RECT 0.000000 11.300000 47.200000 11.500000 ;
      RECT 0.000000 10.700000 46.480000 11.300000 ;
      RECT 0.000000 10.500000 47.200000 10.700000 ;
      RECT 0.000000 9.900000 46.480000 10.500000 ;
      RECT 0.000000 9.700000 47.200000 9.900000 ;
      RECT 0.000000 9.100000 46.480000 9.700000 ;
      RECT 0.000000 8.900000 47.200000 9.100000 ;
      RECT 0.000000 8.300000 46.480000 8.900000 ;
      RECT 0.000000 8.100000 47.200000 8.300000 ;
      RECT 0.000000 7.500000 46.480000 8.100000 ;
      RECT 0.000000 7.300000 47.200000 7.500000 ;
      RECT 0.000000 6.700000 46.480000 7.300000 ;
      RECT 0.000000 6.100000 47.200000 6.700000 ;
      RECT 0.000000 5.500000 46.480000 6.100000 ;
      RECT 0.000000 5.300000 47.200000 5.500000 ;
      RECT 0.000000 4.700000 46.480000 5.300000 ;
      RECT 0.000000 4.500000 47.200000 4.700000 ;
      RECT 0.000000 3.900000 46.480000 4.500000 ;
      RECT 0.000000 3.700000 47.200000 3.900000 ;
      RECT 0.000000 3.100000 46.480000 3.700000 ;
      RECT 0.000000 2.900000 47.200000 3.100000 ;
      RECT 0.000000 2.300000 46.480000 2.900000 ;
      RECT 0.000000 2.100000 47.200000 2.300000 ;
      RECT 0.000000 1.500000 46.480000 2.100000 ;
      RECT 0.000000 1.300000 47.200000 1.500000 ;
      RECT 0.000000 0.700000 46.480000 1.300000 ;
      RECT 0.000000 0.500000 47.200000 0.700000 ;
      RECT 0.000000 0.000000 46.480000 0.500000 ;
    LAYER metal4 ;
      RECT 24.500000 67.280000 47.200000 68.000000 ;
      RECT 20.500000 67.280000 23.900000 68.000000 ;
      RECT 0.000000 67.280000 19.900000 68.000000 ;
      RECT 0.000000 0.720000 47.200000 67.280000 ;
      RECT 24.100000 0.000000 47.200000 0.720000 ;
      RECT 0.000000 0.000000 23.500000 0.720000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 47.200000 68.000000 ;
  END
END BATCHARGERctr

END LIBRARY
