##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Mon Jan 16 11:25:24 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERcore
  CLASS BLOCK ;
  SIZE 640.000000 BY 470.000000 ;
  FOREIGN BATCHARGERcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN iforcedbat
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 296.000000 469.480000 374.000000 470.000000 ;
    END
  END iforcedbat
  PIN vsensbat
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 228.800000 0.000000 230.800000 0.520000 ;
    END
  END vsensbat
  PIN vin
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 285.200000 0.520000 335.200000 ;
    END
  END vin
  PIN vbattemp
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 232.800000 0.000000 234.800000 0.520000 ;
    END
  END vbattemp
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 312.000000 0.000000 312.400000 0.520000 ;
    END
  END en
  PIN sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 316.000000 0.000000 316.400000 0.520000 ;
    END
  END sel[3]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 320.000000 0.000000 320.400000 0.520000 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 324.000000 0.000000 324.400000 0.520000 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 328.000000 0.000000 328.400000 0.520000 ;
    END
  END sel[0]
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 639.480000 24.000000 640.000000 26.000000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 639.480000 29.200000 640.000000 31.200000 ;
    END
  END dgnd
  PIN pgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 159.200000 0.520000 161.200000 ;
    END
  END pgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
    LAYER metal3 ;
      RECT 0.000000 335.480000 640.000000 470.000000 ;
      RECT 0.800000 284.920000 640.000000 335.480000 ;
      RECT 0.000000 161.480000 640.000000 284.920000 ;
      RECT 0.800000 158.920000 640.000000 161.480000 ;
      RECT 0.000000 31.480000 640.000000 158.920000 ;
      RECT 0.000000 28.920000 639.200000 31.480000 ;
      RECT 0.000000 26.280000 640.000000 28.920000 ;
      RECT 0.000000 23.720000 639.200000 26.280000 ;
      RECT 0.000000 0.000000 640.000000 23.720000 ;
    LAYER metal4 ;
      RECT 374.280000 469.200000 640.000000 470.000000 ;
      RECT 0.000000 469.200000 295.720000 470.000000 ;
      RECT 0.000000 0.800000 640.000000 469.200000 ;
      RECT 235.080000 0.720000 640.000000 0.800000 ;
      RECT 328.600000 0.000000 640.000000 0.720000 ;
      RECT 324.600000 0.000000 327.800000 0.720000 ;
      RECT 320.600000 0.000000 323.800000 0.720000 ;
      RECT 316.600000 0.000000 319.800000 0.720000 ;
      RECT 312.600000 0.000000 315.800000 0.720000 ;
      RECT 235.080000 0.000000 311.800000 0.720000 ;
      RECT 231.080000 0.000000 232.520000 0.800000 ;
      RECT 0.000000 0.000000 228.520000 0.800000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 640.000000 470.000000 ;
  END
END BATCHARGERcore

END LIBRARY
